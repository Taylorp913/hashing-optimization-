`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:51:58 02/10/2016 
// Design Name: 
// Module Name:    md5_top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
 module md5_top(port, Clk);

output reg port;
input Clk;

wire [31:0] A0, B0, C0, D0, A, B, C, D, Afin, Bfin, Cfin, Dfin, Atar, Btar, Ctar, Dtar,
		A11, B11, C11, D11, A12, B12, C12, D12, //Round 1 Wires
		A13, B13, C13, D13, A14, B14, C14, D14,
		A15, B15, C15, D15, A16, B16, C16, D16,
		A17, B17, C17, D17, A18, B18, C18, D18,
		A19, B19, C19, D19, A110, B110, C110, D110,
		A111, B111, C111, D111, A112, B112, C112, D112,
		A113, B113, C113, D113, A114, B114, C114, D114,
		A115, B115, C115, D115, A116, B116, C116, D116,
		A21, B21, C21, D21, A22, B22, C22, D22, //Round2 Wires
		A23, B23, C23, D23, A24, B24, C24, D24,
		A25, B25, C25, D25, A26, B26, C26, D26,
		A27, B27, C27, D27, A28, B28, C28, D28,
		A29, B29, C29, D29, A210, B210, C210, D210,
		A211, B211, C211, D211, A212, B212, C212, D212,
		A213, B213, C213, D213, A214, B214, C214, D214,
		A215, B215, C215, D215, A216, B216, C216, D216,
		A31, B31, C31, D31, A32, B32, C32, D32, //Round3 Wires
		A33, B33, C33, D33, A34, B34, C34, D34,
		A35, B35, C35, D35, A36, B36, C36, D36,
		A37, B37, C37, D37, A38, B38, C38, D38,
		A39, B39, C39, D39, A310, B310, C310, D310,
		A311, B311, C311, D311, A312, B312, C312, D312,
		A313, B313, C313, D313, A314, B314, C314, D314,
		A315, B315, C315, D315, A316, B316, C316, D316,
		A41, B41, C41, D41, A42, B42, C42, D42, //Round4 Wires
		A43, B43, C43, D43, A44, B44, C44, D44,
		A45, B45, C45, D45, A46, B46, C46, D46,
		A47, B47, C47, D47, A48, B48, C48, D48,
		A49, B49, C49, D49, A410, B410, C410, D410,
		A411, B411, C411, D411, A412, B412, C412, D412,
		A413, B413, C413, D413, A414, B414, C414, D414,
		A415, B415, C415, D415, A416, B416, C416, D416;
		
		
		
		
		
wire [511:0] X;
wire co;

reg [4:0] K0, K1, K2, K3, K4, K5, K6, K7, K8, K9, K10, K11, K12, K13, K14, K15, K16, K17, K18, K19, K20,
				K21, K22, K23, K24, K25, K26, K27, K28, K29, K30, K31, K32, K33, K34, K35, K36, K37, K38, K39, K40,
				K41, K42, K43, K44, K45, K46, K47, K48, K49, K50,K51, K52, K53, K54, K55, K56, K57, K58, K59, K60, K61, K62, K63, K64;
				
reg [6:0] iter = 0;
reg [6:0] next = 0;
reg [6:0] count = 0;
				
				
				

assign A0[31:0] = 32'h67452301;
assign B0[31:0] = 32'hefcdab89;
assign C0[31:0] = 32'h98badcfe;
assign D0[31:0] = 32'h10325476;

assign A[31:0] = A0[31:0];
assign B[31:0] = B0[31:0];
assign C[31:0] = C0[31:0];
assign D[31:0] = D0[31:0];

assign Atar[31:0] = 32'h0e7a4e0b;
assign Btar[31:0] = 32'hd34ae85f;
assign Ctar[31:0] = 32'h5bf9b55f;
assign Dtar[31:0] = 32'h79acee9c;



//Message for 'aaaaaa'
assign	X[31:0] = 32'h61616161; 	//0
assign	X[63:32] = 32'h00806161; 	//1
assign	X[95:64] = 32'h00000000;	//2
assign	X[127:96] = 32'h00000000;	//3
assign	X[159:128] = 32'h00000000;	//4
assign	X[191:160] = 32'h00000000;	//5
assign	X[223:192] = 32'h00000000;	//6
assign	X[255:224] = 32'h00000000;	//7
assign	X[287:256] = 32'h00000000;	//8
assign	X[319:288] = 32'h00000000;	//9
assign	X[351:320] = 32'h00000000;	//10
assign	X[383:352] = 32'h00000000;	//11
assign	X[415:384] = 32'h00000000;	//12
assign	X[447:416] = 32'h00000000;	//13
assign	X[479:448] = 32'h00000030;	//14
assign	X[511:480] = 32'h00000000;	//15

//Shift array (To make the code more "time dependent")

always@(*) begin
	next[6:0] = iter[6:0] + 1;
	end
	
always@(posedge Clk) begin
		iter[6:0] = next[6:0];
end


always@(*) 
begin
	case(iter[6:0])
	0: K0 = 7;
	1: K1 = 12;
	2: K2 = 17;
	3: K3 = 22;
	4: K4 = 7;
	5: K5 = 12;
	6: K6 = 17;
	7: K7 = 22;
	8: K8 = 7;
	9: K9 = 12;
	10: K10 = 17;
	11: K11 = 22;
	12: K12 = 7;
	13: K13 = 12;
	14: K14 = 17;
	15: K15 = 22; //End of Round 1
	16: K16 = 5;
	17: K17 = 9;
	18: K18 = 14;
	19: K19 = 20;
	20: K20 = 5;
	21: K21 = 9;
	22: K22 = 14;
	23: K23 = 20;
	24: K24 = 5;
	25: K25 = 9;
	26: K26 = 14;
	27: K27 = 20;
	28: K28 = 5;
	29: K29 = 9;
	30: K30 = 14;
	31: K31 = 20; // End of Round 2
	32: K32 = 4;
	33: K33 = 11;
	34: K34 = 16;
	35: K35 = 23;
	36: K36 = 4;
	37: K37 = 11;
	38: K38 = 16;
	39: K39 = 23;
	40: K40 = 4;
	41: K41 = 11;
	42: K42 = 16;
	43: K43 = 23;
	44: K44 = 4;
	45: K45 = 11;
	46: K46 = 16;
	47: K47 = 23; //End of Round 3
	48: K48 = 6;
	49: K49 = 10;
	50: K50 = 15;
	51: K51 = 21;
	52: K52 = 6;
	53: K53 = 10;
	54: K54 = 15;
	55: K55 = 21;
	56: K56 = 6;
	57: K57 = 10;
	58: K58 = 15;
	59: K59 = 21;
	60: K60 = 6;
	61: K61 = 10;
	62: K62 = 15;
	63: K63 = 21;
	default:$display("ERROR IN CASE STATEMENT");
	endcase

end

//Round 1 Function

round1 R11(A11[31:0], B11[31:0], C11[31:0], D11[31:0], A[31:0], B[31:0], C[31:0], D[31:0], X[31:0],  K0, 32'hd76aa478);
round1 R12(A12[31:0], B12[31:0], C12[31:0], D12[31:0], A11[31:0], B11[31:0], C11[31:0], D11[31:0], X[63:32], K1, 32'he8c7b756);
round1 R13(A13[31:0], B13[31:0], C13[31:0], D13[31:0], A12[31:0], B12[31:0], C12[31:0], D12[31:0], X[95:64], K2, 32'h242070db);
round1 R14(A14[31:0], B14[31:0], C14[31:0], D14[31:0], A13[31:0], B13[31:0], C13[31:0], D13[31:0], X[127:96], K3, 32'hc1bdceee);
    
round1 R15(A15[31:0], B15[31:0], C15[31:0], D15[31:0], A14[31:0], B14[31:0], C14[31:0], D14[31:0], X[159:128],  K4, 32'hf57c0faf);
round1 R16(A16[31:0], B16[31:0], C16[31:0], D16[31:0], A15[31:0], B15[31:0], C15[31:0], D15[31:0], X[191:160], K5, 32'h4787c62a);
round1 R17(A17[31:0], B17[31:0], C17[31:0], D17[31:0], A16[31:0], B16[31:0], C16[31:0], D16[31:0], X[223:192], K6, 32'ha8304613);
round1 R18(A18[31:0], B18[31:0], C18[31:0], D18[31:0], A17[31:0], B17[31:0], C17[31:0], D17[31:0], X[255:224], K7, 32'hfd469501);

round1 R19(A19[31:0],  B19[31:0], C19[31:0], D19[31:0], A18[31:0], B18[31:0], C18[31:0], D18[31:0], X[287:256],  K8, 32'h698098d8);
round1 R110(A110[31:0], B110[31:0], C110[31:0], D110[31:0], A19[31:0], B19[31:0], C19[31:0], D19[31:0], X[319:288], K9, 32'h8b44f7af);
round1 R111(A111[31:0], B111[31:0], C111[31:0], D111[31:0], A110[31:0], B110[31:0], C110[31:0], D110[31:0], X[351:320], K10, 32'hffff5bb1);
round1 R112(A112[31:0], B112[31:0], C112[31:0], D112[31:0], A111[31:0], B111[31:0], C111[31:0], D111[31:0], X[383:352], K11, 32'h895cd7be);
   
round1 R113(A113[31:0], B113[31:0], C113[31:0], D113[31:0], A112[31:0], B112[31:0], C112[31:0], D112[31:0], X[415:384], K12, 32'h6b901122);
round1 R114(A114[31:0], B114[31:0], C114[31:0], D114[31:0], A113[31:0], B113[31:0], C113[31:0], D113[31:0], X[447:416],K13, 32'hfd987193);
round1 R115(A115[31:0], B115[31:0], C115[31:0], D115[31:0], A114[31:0], B114[31:0], C114[31:0], D114[31:0], X[479:448],K14, 32'ha679438e);
round1 R116(A116[31:0], B116[31:0], C116[31:0], D116[31:0], A115[31:0], B115[31:0], C115[31:0], D115[31:0], X[511:480],K15, 32'h49b40821);

 
//Round 2 Functions
round2 R21(A21[31:0], B21[31:0], C21[31:0], D21[31:0], A116[31:0], B116[31:0], C116[31:0], D116[31:0], X[63:32],    K16, 32'hf61e2562);
round2 R22(A22[31:0], B22[31:0], C22[31:0], D22[31:0], A21[31:0], B21[31:0], C21[31:0], D21[31:0], X[223:192],      K17, 32'hc040b340);
round2 R23(A23[31:0], B23[31:0], C23[31:0], D23[31:0], A22[31:0], B22[31:0], C22[31:0], D22[31:0], X[383:352],     K18, 32'h265e5a51);
round2 R24(A24[31:0], B24[31:0], C24[31:0], D24[31:0], A23[31:0], B23[31:0], C23[31:0], D23[31:0], X[31:0],        K19, 32'he9b6c7aa);
 
round2 R25(A25[31:0], B25[31:0], C25[31:0], D25[31:0], A24[31:0], B24[31:0], C24[31:0], D24[31:0], X[191:160],      K20, 32'hd62f105d);
round2 R26(A26[31:0], B26[31:0], C26[31:0], D26[31:0], A25[31:0], B25[31:0], C25[31:0], D25[31:0], X[351:320],      K21, 32'h02441453);
round2 R27(A27[31:0], B27[31:0], C27[31:0], D27[31:0], A26[31:0], B26[31:0], C26[31:0], D26[31:0], X[511:480],     K22, 32'hd8a1e681);
round2 R28(A28[31:0], B28[31:0], C28[31:0], D28[31:0], A27[31:0], B27[31:0], C27[31:0], D27[31:0], X[159:128],     K23, 32'he7d3fbc8);
    
round2 R29(A29[31:0], B29[31:0], C29[31:0], D29[31:0], A28[31:0], B28[31:0], C28[31:0], D28[31:0], X[319:288],          K24, 32'h21e1cde6);
round2 R210(A210[31:0], B210[31:0], C210[31:0], D210[31:0], A29[31:0], B29[31:0], C29[31:0], D29[31:0], X[479:448],     K25, 32'hc33707d6);
round2 R211(A211[31:0], B211[31:0], C211[31:0], D211[31:0], A210[31:0], B210[31:0], C210[31:0], D210[31:0], X[127:96], K26, 32'hf4d50d87);
round2 R212(A212[31:0], B212[31:0], C212[31:0], D212[31:0], A211[31:0], B211[31:0], C211[31:0], D211[31:0], X[287:256], K27, 32'h455a14ed);
    
round2 R213(A213[31:0], B213[31:0], C213[31:0], D213[31:0], A212[31:0], B212[31:0], C212[31:0], D212[31:0], X[447:416],  K28, 32'ha9e3e905);
round2 R214(A214[31:0], B214[31:0], C214[31:0], D214[31:0], A213[31:0], B213[31:0], C213[31:0], D213[31:0], X[95:64],    K29, 32'hfcefa3f8);
round2 R215(A215[31:0], B215[31:0], C215[31:0], D215[31:0], A214[31:0], B214[31:0], C214[31:0], D214[31:0], X[255:224], K30, 32'h676f02d9);
round2 R216(A216[31:0], B216[31:0], C216[31:0], D216[31:0], A215[31:0], B215[31:0], C215[31:0], D215[31:0], X[415:384], K31, 32'h8d2a4c8a);
    
    
//Round 3 Functions 
round3 R31(A31[31:0], B31[31:0], C31[31:0], D31[31:0], A216[31:0], B216[31:0], C216[31:0], D216[31:0], X[191:160],  K32, 32'hfffa3942);
round3 R32(A32[31:0], B32[31:0], C32[31:0], D32[31:0], A31[31:0], B31[31:0], C31[31:0], D31[31:0], X[287:256], K33, 32'h8771f681);
round3 R33(A33[31:0], B33[31:0], C33[31:0], D33[31:0], A32[31:0], B32[31:0], C32[31:0], D32[31:0], X[383:352], K34, 32'h6d9d6122);
round3 R34(A34[31:0], B34[31:0], C34[31:0], D34[31:0], A33[31:0], B33[31:0], C33[31:0], D33[31:0], X[479:448], K35, 32'hfde5380c);
   
round3 R35(A35[31:0], B35[31:0], C35[31:0], D35[31:0], A34[31:0], B34[31:0], C34[31:0], D34[31:0], X[63:32],  K36, 32'ha4beea44);
round3 R36(A36[31:0], B36[31:0], C36[31:0], D36[31:0], A35[31:0], B35[31:0], C35[31:0], D35[31:0], X[159:128], K37, 32'h4bdecfa9);
round3 R37(A37[31:0], B37[31:0], C37[31:0], D37[31:0], A36[31:0], B36[31:0], C36[31:0], D36[31:0], X[255:224], K38, 32'hf6bb4b60);
round3 R38(A38[31:0], B38[31:0], C38[31:0], D38[31:0], A37[31:0], B37[31:0], C37[31:0], D37[31:0], X[351:320], K39, 32'hbebfbc70);
    
round3 R39(A39[31:0], B39[31:0], C39[31:0], D39[31:0], A38[31:0], B38[31:0], C38[31:0], D38[31:0], X[447:416], K40, 32'h289b7ec6);
round3 R310(A310[31:0], B310[31:0], C310[31:0], D310[31:0], A39[31:0], B39[31:0], C39[31:0], D39[31:0],X[31:0], K41, 32'heaa127fa);
round3 R311(A311[31:0], B311[31:0], C311[31:0], D311[31:0], A310[31:0], B310[31:0], C310[31:0], D310[31:0], X[127:96], K42, 32'hd4ef3085);
round3 R312(A312[31:0], B312[31:0], C312[31:0], D312[31:0], A311[31:0], B311[31:0], C311[31:0], D311[31:0], X[223:192], K43, 32'h04881d05);
    
round3 R313(A313[31:0], B313[31:0], C313[31:0], D313[31:0], A312[31:0], B312[31:0], C312[31:0], D312[31:0], X[319:288],  K44, 32'hd9d4d039);
round3 R314(A314[31:0], B314[31:0], C314[31:0], D314[31:0], A313[31:0], B313[31:0], C313[31:0], D313[31:0], X[415:384], K45, 32'he6db99e5);
round3 R315(A315[31:0], B315[31:0], C315[31:0], D315[31:0], A314[31:0], B314[31:0], C314[31:0], D314[31:0], X[511:480], K46, 32'h1fa27cf8);
round3 R316(A316[31:0], B316[31:0], C316[31:0], D316[31:0], A315[31:0], B315[31:0], C315[31:0], D315[31:0], X[95:64],  K47, 32'hc4ac5665);
    
    
 
round4 R41(A41[31:0], B41[31:0], C41[31:0], D41[31:0], A316[31:0], B316[31:0], C316[31:0], D316[31:0], X[31:0],  K48, 32'hf4292244);
round4 R42(A42[31:0], B42[31:0], C42[31:0], D42[31:0], A41[31:0], B41[31:0], C41[31:0], D41[31:0], X[255:224], K49, 32'h432aff97);
round4 R43(A43[31:0], B43[31:0], C43[31:0], D43[31:0], A42[31:0], B42[31:0], C42[31:0], D42[31:0], X[479:448], K50, 32'hab9423a7);
round4 R44(A44[31:0], B44[31:0], C44[31:0], D44[31:0], A43[31:0], B43[31:0], C43[31:0], D43[31:0], X[191:160], K51, 32'hfc93a039);
    
round4 R45(A45[31:0], B45[31:0], C45[31:0], D45[31:0], A44[31:0], B44[31:0], C44[31:0], D44[31:0], X[415:384], K52, 32'h655b59c3);
round4 R46(A46[31:0], B46[31:0], C46[31:0], D46[31:0], A45[31:0], B45[31:0], C45[31:0], D45[31:0], X[127:96], K53, 32'h8f0ccc92);
round4 R47(A47[31:0], B47[31:0], C47[31:0], D47[31:0], A46[31:0], B46[31:0], C46[31:0], D46[31:0], X[351:320],K54, 32'hffeff47d);
round4 R48(A48[31:0], B48[31:0], C48[31:0], D48[31:0], A47[31:0], B47[31:0], C47[31:0], D47[31:0], X[63:32], K55, 32'h85845dd1);
    
round4 R49(A49[31:0], B49[31:0], C49[31:0], D49[31:0], A48[31:0], B48[31:0], C48[31:0], D48[31:0], X[287:256],  K56, 32'h6fa87e4f);
round4 R410(A410[31:0], B410[31:0], C410[31:0], D410[31:0], A49[31:0], B49[31:0], C49[31:0], D49[31:0], X[511:480], K57, 32'hfe2ce6e0);
round4 R411(A411[31:0], B411[31:0], C411[31:0], D411[31:0], A410[31:0], B410[31:0], C410[31:0], D410[31:0], X[223:192], K58, 32'ha3014314);
round4 R412(A412[31:0], B412[31:0], C412[31:0], D412[31:0], A411[31:0], B411[31:0], C411[31:0], D411[31:0], X[447:416], K59, 32'h4e0811a1);
    
round4 R413(A413[31:0], B413[31:0], C413[31:0], D413[31:0], A412[31:0], B412[31:0], C412[31:0], D412[31:0], X[159:128],  K60, 32'hf7537e82);
round4 R414(A414[31:0], B414[31:0], C414[31:0], D414[31:0], A413[31:0], B413[31:0], C413[31:0], D413[31:0], X[383:352], K61, 32'hbd3af235);
round4 R415(A415[31:0], B415[31:0], C415[31:0], D415[31:0], A414[31:0], B414[31:0], C414[31:0], D414[31:0], X[95:64], K62, 32'h2ad7d2bb);
round4 R416(A416[31:0], B416[31:0], C416[31:0], D416[31:0], A415[31:0], B415[31:0], C415[31:0], D415[31:0], X[319:288], K63, 32'heb86d391);
	 

assign Afin[31:0] = A416[31:0] + A0[31:0];
assign Bfin[31:0] = B416[31:0] + B0[31:0];
assign Cfin[31:0] = C416[31:0] + C0[31:0];
assign Dfin[31:0] = D416[31:0] + D0[31:0];

	 
always@(posedge Clk) begin
	if(Afin[31:0] == Atar[31:0] && Bfin[31:0] == Btar[31:0] && Cfin[31:0] == Ctar[31:0] && Dfin[31:0] == Dtar[31:0]) begin
	port <= 1;
	end
end
	


endmodule
